`ifndef __GLOSSY_VH__
`define __GLOSSY_VH__

`define GLOSSY_RXTX_ADDR_FRM_START       7'h00
`define GLOSSY_RXTX_ADDR_FRM_LEN         7'h00
`define GLOSSY_RXTX_ADDR_RL_CNT          7'h01
`define GLOSSY_RXTX_ADDR_DATA_START      7'h02

`endif // __GLOSSY_VH__