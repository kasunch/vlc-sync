`ifndef __TX_VH__
`define __TX_VH__

`define TX_EVENT_NONE           3'd0
`define TX_EVENT_STARTED        3'd1
`define TX_EVENT_PREAMBLE       3'd2
`define TX_EVENT_SFD            3'd3
`define TX_EVENT_PHR            3'h4
`define TX_EVENT_BYTE           3'h5
`define TX_EVENT_END            3'h6

`endif // __TX_VH__
