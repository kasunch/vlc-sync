`ifndef __RX_TB_VH__
`define __RX_TB_VH__

`define RX_INPUT_DATA_SIZE  10000

`endif // __RX_TB_VH__