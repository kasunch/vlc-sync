`ifndef __SYM_COMMON_VH__
`define __SYM_COMMON_VH__

//`define SYM_ENC_DEC_PREAMBLE            8'hAA
`define SYM_ENC_DEC_PREAMBLE            8'h00   
`define SYM_ENC_DEC_SFD                 8'h11

`define SYM_ENC_DEC_PREAMBLE_SIZE       8
`define SYM_ENC_DEC_SFD_SIZE            8      
`define SYM_ENC_DEC_PHR_SIZE            8      
`define SYM_ENC_DEC_FCS_SIZE            16

`endif // __SYM_COMMON_VH__