`ifndef __UART_CFG_VH__
`define __UART_CFG_VH__

`define CLKS_PER_BIT_115200   347

`endif // __UART_CFG_VH__