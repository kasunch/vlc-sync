module schmidl_cox_preamble(clk, reset, i_r_addr, o_data);
    input clk;
    input reset;
    input [7:0] i_r_addr;
    output reg [9:0] o_data;

    always @(posedge clk) begin
        case (i_r_addr)
            8'h000 : o_data <= 10'h200;
            8'h001 : o_data <= 10'h1E2;
            8'h002 : o_data <= 10'h2E3;
            8'h003 : o_data <= 10'h1D9;
            8'h004 : o_data <= 10'h1CF;
            8'h005 : o_data <= 10'h218;
            8'h006 : o_data <= 10'h140;
            8'h007 : o_data <= 10'h0EC;
            8'h008 : o_data <= 10'h213;
            8'h009 : o_data <= 10'h1BF;
            8'h00A : o_data <= 10'h2B1;
            8'h00B : o_data <= 10'h0EA;
            8'h00C : o_data <= 10'h2ED;
            8'h00D : o_data <= 10'h148;
            8'h00E : o_data <= 10'h15D;
            8'h00F : o_data <= 10'h01A;
            8'h010 : o_data <= 10'h128;
            8'h011 : o_data <= 10'h1DC;
            8'h012 : o_data <= 10'h2F2;
            8'h013 : o_data <= 10'h237;
            8'h014 : o_data <= 10'h1C3;
            8'h015 : o_data <= 10'h27F;
            8'h016 : o_data <= 10'h06A;
            8'h017 : o_data <= 10'h1FB;
            8'h018 : o_data <= 10'h3A8;
            8'h019 : o_data <= 10'h1D4;
            8'h01A : o_data <= 10'h217;
            8'h01B : o_data <= 10'h232;
            8'h01C : o_data <= 10'h17F;
            8'h01D : o_data <= 10'h0BA;
            8'h01E : o_data <= 10'h17A;
            8'h01F : o_data <= 10'h205;
            8'h020 : o_data <= 10'h17A;
            8'h021 : o_data <= 10'h0BA;
            8'h022 : o_data <= 10'h17F;
            8'h023 : o_data <= 10'h232;
            8'h024 : o_data <= 10'h217;
            8'h025 : o_data <= 10'h1D4;
            8'h026 : o_data <= 10'h3A8;
            8'h027 : o_data <= 10'h1FB;
            8'h028 : o_data <= 10'h06A;
            8'h029 : o_data <= 10'h27F;
            8'h02A : o_data <= 10'h1C3;
            8'h02B : o_data <= 10'h237;
            8'h02C : o_data <= 10'h2F2;
            8'h02D : o_data <= 10'h1DC;
            8'h02E : o_data <= 10'h128;
            8'h02F : o_data <= 10'h01A;
            8'h030 : o_data <= 10'h15D;
            8'h031 : o_data <= 10'h148;
            8'h032 : o_data <= 10'h2ED;
            8'h033 : o_data <= 10'h0EA;
            8'h034 : o_data <= 10'h2B1;
            8'h035 : o_data <= 10'h1BF;
            8'h036 : o_data <= 10'h213;
            8'h037 : o_data <= 10'h0EC;
            8'h038 : o_data <= 10'h140;
            8'h039 : o_data <= 10'h218;
            8'h03A : o_data <= 10'h1CF;
            8'h03B : o_data <= 10'h1D9;
            8'h03C : o_data <= 10'h2E3;
            8'h03D : o_data <= 10'h1E2;
            8'h03E : o_data <= 10'h200;
            8'h03F : o_data <= 10'h200;
            8'h040 : o_data <= 10'h200;
            8'h041 : o_data <= 10'h1E2;
            8'h042 : o_data <= 10'h2E3;
            8'h043 : o_data <= 10'h1D9;
            8'h044 : o_data <= 10'h1CF;
            8'h045 : o_data <= 10'h218;
            8'h046 : o_data <= 10'h140;
            8'h047 : o_data <= 10'h0EC;
            8'h048 : o_data <= 10'h213;
            8'h049 : o_data <= 10'h1BF;
            8'h04A : o_data <= 10'h2B1;
            8'h04B : o_data <= 10'h0EA;
            8'h04C : o_data <= 10'h2ED;
            8'h04D : o_data <= 10'h148;
            8'h04E : o_data <= 10'h15D;
            8'h04F : o_data <= 10'h01A;
            8'h050 : o_data <= 10'h128;
            8'h051 : o_data <= 10'h1DC;
            8'h052 : o_data <= 10'h2F2;
            8'h053 : o_data <= 10'h237;
            8'h054 : o_data <= 10'h1C3;
            8'h055 : o_data <= 10'h27F;
            8'h056 : o_data <= 10'h06A;
            8'h057 : o_data <= 10'h1FB;
            8'h058 : o_data <= 10'h3A8;
            8'h059 : o_data <= 10'h1D4;
            8'h05A : o_data <= 10'h217;
            8'h05B : o_data <= 10'h232;
            8'h05C : o_data <= 10'h17F;
            8'h05D : o_data <= 10'h0BA;
            8'h05E : o_data <= 10'h17A;
            8'h05F : o_data <= 10'h205;
            8'h060 : o_data <= 10'h17A;
            8'h061 : o_data <= 10'h0BA;
            8'h062 : o_data <= 10'h17F;
            8'h063 : o_data <= 10'h232;
            8'h064 : o_data <= 10'h217;
            8'h065 : o_data <= 10'h1D4;
            8'h066 : o_data <= 10'h3A8;
            8'h067 : o_data <= 10'h1FB;
            8'h068 : o_data <= 10'h06A;
            8'h069 : o_data <= 10'h27F;
            8'h06A : o_data <= 10'h1C3;
            8'h06B : o_data <= 10'h237;
            8'h06C : o_data <= 10'h2F2;
            8'h06D : o_data <= 10'h1DC;
            8'h06E : o_data <= 10'h128;
            8'h06F : o_data <= 10'h01A;
            8'h070 : o_data <= 10'h15D;
            8'h071 : o_data <= 10'h148;
            8'h072 : o_data <= 10'h2ED;
            8'h073 : o_data <= 10'h0EA;
            8'h074 : o_data <= 10'h2B1;
            8'h075 : o_data <= 10'h1BF;
            8'h076 : o_data <= 10'h213;
            8'h077 : o_data <= 10'h0EC;
            8'h078 : o_data <= 10'h140;
            8'h079 : o_data <= 10'h218;
            8'h07A : o_data <= 10'h1CF;
            8'h07B : o_data <= 10'h1D9;
            8'h07C : o_data <= 10'h2E3;
            8'h07D : o_data <= 10'h1E2;
            8'h07E : o_data <= 10'h200;
            8'h07F : o_data <= 10'h200;
            default: o_data <= 0;
        endcase
    end
endmodule
