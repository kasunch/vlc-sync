`ifndef __RX_VH__
`define __RX_VH__

`define RX_EVENT_NONE           3'd0
`define RX_EVENT_PREAMBLE       3'd1
`define RX_EVENT_SFD            3'd2
`define RX_EVENT_PHR            3'h3
`define RX_EVENT_BYTE           3'h4
`define RX_EVENT_END            3'h5

`endif // __RX_VH__
