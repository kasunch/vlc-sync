`ifndef __SYM_ENC_VH__
`define __SYM_ENC_VH__

`define SYM_ENC_EV_NONE        3'd0
`define SYM_ENC_EV_STARTED     3'd1
`define SYM_ENC_EV_PREAMBLE    3'd2
`define SYM_ENC_EV_SFD         3'd3
`define SYM_ENC_EV_PHR         3'd4
`define SYM_ENC_EV_BYTE        3'd5
`define SYM_ENC_EV_COMPLETE    3'd6

`endif // __SYM_ENC_VH__
